hi this is disturbing
