hey there this is another test
